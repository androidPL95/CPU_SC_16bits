library verilog;
use verilog.vl_types.all;
entity typedefs is
end typedefs;
