library verilog;
use verilog.vl_types.all;
entity SingleCycle_Top_tb is
end SingleCycle_Top_tb;
